module decoder();
/*	assign iv = d[23:8];
	assign as = d[7]; ms, mwe, rwe,
	assign aaddr = d[6:5];
	assign baddr = d[4:3];
	assign op = d[2];
	assign oaddr = d[1:0];
*/
endmodule