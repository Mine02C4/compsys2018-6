module imem(addr, d);
	input [7:0] addr;
	output [23:0] d;
	reg [23:0] d;
//  a[2], b[2], op[1], o[2]
	always @(*) begin
		case (addr)
	8'h00: d = 24'b0000000000000001_1_00_00_1_00;
	8'h01: d = 24'b0000000000000001_1_00_00_1_01;
	8'h02: d = 24'b0000000000000000_0_00_01_1_10;
	8'h03: d = 24'b0000000000000000_0_01_00_0_00;
	8'h04: d = 24'b0000000000000000_0_10_00_0_01;
	8'h05: d = 24'b0000000000000000_0_00_01_1_10;
	8'h06: d = 24'b0000000000000000_0_01_00_0_00;
	8'h07: d = 24'b0000000000000000_0_10_00_0_01;
	8'h08: d = 24'b0000000000000000_0_00_01_1_10;
	8'h09: d = 24'b0000000000000000_0_01_00_0_00;
	8'h0a: d = 24'b0000000000000000_0_10_00_0_01;
	8'h0b: d = 24'b0000000000000000_0_00_01_1_10;
	8'h0c: d = 24'b0000000000000000_0_01_00_0_00;
	8'h0d: d = 24'b0000000000000000_0_10_00_0_01;
	8'h0e: d = 24'b0000000000000000_0_00_01_1_10;
	8'h0f: d = 24'b0000000000000000_0_01_00_0_00;
	8'h10: d = 24'b0000000000000000_0_10_00_0_01;
	8'h11: d = 24'b0000000000000000_0_00_01_1_10;
	8'h12: d = 24'b0000000000000000_0_01_00_0_00;
	8'h13: d = 24'b0000000000000000_0_10_00_0_01;
	8'h14: d = 24'b0000000000000000_0_00_01_1_10;
	8'h15: d = 24'b0000000000000000_0_01_00_0_00;
	8'h16: d = 24'b0000000000000000_0_10_00_0_01;
		endcase
	end
endmodule
